// Sample source; could use external/lib.v via symlink
module main;
endmodule
