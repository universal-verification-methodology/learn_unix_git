// Sample source for clean_build example
module main;
endmodule
