// Sample testbench for makefile_basics example
module test_main;
endmodule
