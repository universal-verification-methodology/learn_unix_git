// Sample for Module 5 find_grep example.
// Does not contain CLOCK_SIGNAL.
module util (input a, output b);
  assign b = ~a;
endmodule
