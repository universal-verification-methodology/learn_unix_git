// sample design for wildcard example
module design;
endmodule
