// Sample testbench for clean_build example
module test_main;
endmodule
