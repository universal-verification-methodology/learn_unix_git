// Shared library for link_relative example
module lib;
endmodule
