// Sample source for makefile_basics example
module main;
endmodule
